//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Tue Aug 12 00:02:00 2025
// Version: 2024.2 2024.2.0.13
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// mat
module mat(
    // Inputs
    A,
    B,
    clk,
    rst,
    // Outputs
    C
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  [31:0] A;
input  [31:0] B;
input         clk;
input         rst;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [31:0] C;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   [31:0] A;
wire   [31:0] B;
wire   [31:0] C_net_0;
wire          clk;
wire          rst;
wire   [31:0] C_net_1;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign C_net_1 = C_net_0;
assign C[31:0] = C_net_1;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------matmul
matmul matmul_0(
        // Inputs
        .clk ( clk ),
        .rst ( rst ),
        .A   ( A ),
        .B   ( B ),
        // Outputs
        .C   ( C_net_0 ) 
        );


endmodule
