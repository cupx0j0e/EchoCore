-- This is automatically generated INCLUDE (Verilog)
-- or Package (VHDL) file of Enum FIR const coeffs
-- Model ROM's for PHY_TAPS MAC's.  Images of the ROM's are 
-- depicted below for example of 99-tap filter.           

-- Tap                    Coef set (ROM Addr)               
--        0       1       2    ...    13      14      15    
--  0   c0_0    c0_1    c0_2        c0_13   c0_14   c0_15 
--  1   c1_0    c1_1    c1_2        c1_13   c1_14   c1_15 
--  2   c2_0    c2_1    c2_2        c2_13   c2_14   c2_15 
-- ...  
--  98  c98_0   c98_1   c98_2       c98_13  c98_14  c98_15

-- To comply with G5 lib, the 16 coefs of the same tap are concateneted into 
-- a single vector of width 16*18=288, e.g.:    
--  {c1_15, c1_14, c1_13, c1_12, ..., c1_2, c1_1, c1_0}  

-- Furthermore, the 288-bit vectors are concatenated into a single flattened 
-- vector of 288*PHY_TAPS bits 
LIBRARY ieee; 
  USE IEEE.std_logic_1164.all; 

PACKAGE fir_hilbert_fir_hilbert_0_enumFIR_coefs IS
 type   mem_t is array(2 downto 0) of std_logic_vector(1727 downto 0) ; 
  constant INIT : mem_t := (   
( "000000000011101110" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & 
"000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & 
"000000010000100000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & 
"000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & 
"000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & 
"000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000"
 ),  
( "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & 
"000001000101110011" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & 
"000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & 
"000100110111000110" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & 
"000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & 
"111011001000111010" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000"
 ),  
( "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & 
"111110111010001101" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & 
"000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & 
"111111101111100000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & 
"000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & 
"111111111100010010" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000" & "000000000000000000"
 ) ) ; 
END fir_hilbert_fir_hilbert_0_enumFIR_coefs;
