`timescale 1ps/1ps

module preproc_tb;



endmodule