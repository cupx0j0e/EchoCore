-- This is automatically generated INCLUDE (Verilog) or Package (VHDL) 
-- file of Enum FIR array-style parameters
-- RC parameters
LIBRARY ieee; 
  USE IEEE.std_logic_1164.all; 

PACKAGE COREFIR_PF_C0_COREFIR_PF_C0_0_enum_params IS
  constant RC_MM_BITS      : integer := 8; 
  constant RC_MAX_MAC_ROWS : integer := 20; 
  constant RC_ROWS  : integer := 1; 
  constant FIRST_ROW_SIZE  : integer := 6; 
  constant HIGH_ROW_SIZE  : integer := 6; 
  constant RC_INFO : std_logic_vector(159 DOWNTO 0) := 
"00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000110"; 
  constant RC_RANK : std_logic_vector(159 DOWNTO 0) := 
"00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000001"; 
  constant RC_ADV_DDLY_D : std_logic_vector(159 DOWNTO 0) := 
"00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000"; 
  constant RC_ADV_DDLY_S : std_logic_vector(159 DOWNTO 0) := 
"00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00000000" & "00001001"; 
END COREFIR_PF_C0_COREFIR_PF_C0_0_enum_params;
