module start_pulse_generator (
    input clk,
    input reset,
    output start_pulse
);
    
    assign start_pulse = 1'b1;

endmodule
