//****************************************************************
//Microsemi Corporation Proprietary and Confidential
//Copyright 2014 Microsemi Corporation.  All rights reserved
//
//ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
//ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE 
//APPROVED IN ADVANCE IN WRITING.
//
//Description: CoreCORDIC
//             Parallel architecture. LUT
//
//Rev:
//v4.0 12/2/2014  Porting in TGI framework
//
//SVN Revision Information:
//SVN$Revision:$
//SVN$Date:$
//
//Resolved SARS
//
//
//
//Notes:
//
//****************************************************************
module CORECORDIC_C0_CORECORDIC_C0_0_cROM_par(arctan, rcprGain_fx);
  parameter DP_BITS = 8;
  parameter ITERATION = 0;

  localparam IN_BITS = 48;

  output[DP_BITS-1:0] arctan;
  output[IN_BITS-1:0] rcprGain_fx;
  generate  
    case (ITERATION)  
      0: assign arctan = 48'b000100000000000000000000000000000000000000000000;  //  48'd17592186044416
      1: assign arctan = 48'b000010010111001000000010100011101100111011111010;  //  48'd10385273835258
      2: assign arctan = 48'b000001001111110110011100001011011010111101110010;  //  48'd5487293476722
      3: assign arctan = 48'b000000101000100010001000111010100000111011101111;  //  48'd2785435848431
      4: assign arctan = 48'b000000010100010110000110101000011000011100101100;  //  48'd1398123104044
      5: assign arctan = 48'b000000001010001011101011111100001010110010000010;  //  48'd699743120514
      6: assign arctan = 48'b000000000101000101111011000011110010111000010100;  //  48'd349956943380
      7: assign arctan = 48'b000000000010100010111110001010101000100011101010;  //  48'd174989150442
      8: assign arctan = 48'b000000000001010001011111001010011010001101101000;  //  48'd87495910248
      9: assign arctan = 48'b000000000000101000101111100101110101110110011000;  //  48'd43748122008
     10: assign arctan = 48'b000000000000010100010111110011000000000001001001;  //  48'd21874081865
     11: assign arctan = 48'b000000000000001010001011111001100000101001010100;  //  48'd10937043540
     12: assign arctan = 48'b000000000000000101000101111100110000011001110000;  //  48'd5468522096
     13: assign arctan = 48'b000000000000000010100010111110011000001101100001;  //  48'd2734261089
     14: assign arctan = 48'b000000000000000001010001011111001100000110110101;  //  48'd1367130549
     15: assign arctan = 48'b000000000000000000101000101111100110000011011011;  //  48'd683565275
      default: assign arctan = 48'b000000000000000000101000101111100110000011011011;  //  48'd683565275
    endcase
  endgenerate
  assign rcprGain_fx = 48'd42731626441408; 
endmodule
