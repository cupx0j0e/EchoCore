module basic_input_output_signal
(
input            in_sig,
output           out_sig
);

assign out_sig = in_sig;

endmodule

